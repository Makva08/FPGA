module displ(
	input enable,
	input [3:0] digit,
	output reg [7:0] display);
	
endmodule
